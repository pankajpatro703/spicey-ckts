CMOS 2-input TG NOR
*
*    Copyright 2020 Pankajkumar Patro Licensed under the
*    Educational Community License, Version 2.0 (the "License"); you may
*    not use this file except in compliance with the License. You may
*    obtain a copy of the License at
*    
*    http://www.osedu.org/licenses/ECL-2.0
*
*    Unless required by applicable law or agreed to in writing,
*    software distributed under the License is distributed on an "AS IS"
*    BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express
*    or implied. See the License for the specific language governing
*    permissions and limitations under the License.
*
***************************
* @Author: pankajpatro703 *
*  Released under ECL v2  *
***************************
vdd 1 0 dc    5v
va  a 0 pulse 0v 5v 0ns 10us 10us 2ms 4ms	*input A
vb  b 0 pulse 0v 5v 0ns 10us 10us 4ms 8ms	*input B
*output at node Y
**********
mcn1 n1 a  0  0  nmod w=10u l=2u
mcn2 n2 b  0  0  nmod w=10u l=2u
mtn1 n2 n1 y  0  nmod w=10u l=2u
mtn2 0  a  y  0  nmod w=10u l=2u
mtp1 y  a  n2 1  pmod w=10u l=2u
mtp2 y  n1 0  1  pmod w=10u l=2u
mcp1 n1 a  1  1  pmod w=10u l=2u
mcp2 n2 b  1  1  pmod w=10u l=2u
**********
.model nmod nmos vto=1v  kp=20u
.model pmod pmos vto=-1v kp=20u
.tran 0ns 8ms 10us 100us
.control
run
plot v(y) v(a) v(b)
.endc
.end
