CMOS 2-input Dynamic NOR
*
*    Copyright 2020 Pankajkumar Patro Licensed under the
*    Educational Community License, Version 2.0 (the "License"); you may
*    not use this file except in compliance with the License. You may
*    obtain a copy of the License at
*    
*    http://www.osedu.org/licenses/ECL-2.0
*
*    Unless required by applicable law or agreed to in writing,
*    software distributed under the License is distributed on an "AS IS"
*    BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express
*    or implied. See the License for the specific language governing
*    permissions and limitations under the License.
*
***************************
* @Author: pankajpatro703 *
*  Released under ECL v2  *
***************************
vdd 1 0 dc 5v
va 2 0 pulse 0v 5v 0ns 10us 10us 1ms 2ms  	*input A
vb 3 0 pulse 0v 5v 0ns 10us 10us 2ms 4ms  	*input B
vk 4 0 pulse 0v 5v 0ns 10us 10us 0.9ms 1ms	*clock phi
*output at node 6
**********
mcn1 6 2 5 0 nmod w=10u l=2u
mcn2 6 3 5 0 nmod w=10u l=2u
mkn1 5 4 0 0 nmod w=10u l=2u
mkp1 6 4 1 1 pmod w=10u l=2u
mbp1 6 6 1 1 pmod w=10u l=40u
**********
.model nmod nmos vto=1v kp=20u
.model pmod pmos vto=-1v kp=20u
.tran 0ns 4ms 10us 100us
.control
run
plot v(6) v(2) v(3)
plot v(4)
.endc
.end
