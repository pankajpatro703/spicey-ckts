CMOS 4-to-1 MUX
*
*    Copyright 2020 Pankajkumar Patro Licensed under the
*    Educational Community License, Version 2.0 (the "License"); you may
*    not use this file except in compliance with the License. You may
*    obtain a copy of the License at
*    
*    http://www.osedu.org/licenses/ECL-2.0
*
*    Unless required by applicable law or agreed to in writing,
*    software distributed under the License is distributed on an "AS IS"
*    BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express
*    or implied. See the License for the specific language governing
*    permissions and limitations under the License.
*
***************************
* @Author: pankajpatro703 *
*  Released under ECL v2  *
***************************
vdd  1   0 dc    5v
vwl  wl  0 pulse 5v 0v 0ns 10us 10us 0.5ms 2ms	*input WordLine
vs   sel 0 pulse 0v 5v 0ns 10us 10us 2ms   4ms	*input SelectLine
vbl  bl  0 pulse 5v 0v 0ns 10us 10us 4ms   8ms	*input BitLine
vbl1 bl1 0 pulse 0v 5v 0ns 10us 10us 4ms   8ms	*complement of BitLine
*output at nodes q, q1, c, c1
**********
cb1 c  0 100pF
cb2 c1 0 100pF
**********
mbn1 c  sel bl  0  nmod w=100u l=2u 
mbn2 c1 sel bl1 0  nmod w=100u l=2u 
mcn2 q  q1  0   0  nmod w=10u  l=2u 
mcn1 q1 q   0   0  nmod w=10u  l=2u 
mcc1 C1 wl  q1  0  nmod w=10u  l=2u 
mcc2 C  wl  q   0  nmod w=10u  l=2u 
mvp1 1  0   c   1  pmod w=10u  l=2u 
mvp2 1  0   c1  1  pmod w=10u  l=2u 
mpn1 1  q   q1  1  pmod w=10u  l=2u 
mpn2 1  q1  q   1  pmod w=10u  l=2u 
**********
.model nmod nmos vto=1v  kp=20u
.model pmod pmos vto=-1v kp=20u
.tran 0ns 8ms 10us 100us
.control
run
plot v(bl) v(sel) v(wl)
plot v(q) v(c)
plot v(q1) v(c1)
.endc
.end
