CMOS 2-input NOR
***************************
* @Author: pankajpatro703 *
*  Released under ECL v2  *
***************************
vdd 1 0 dc 5v
va 3 0 pulse 0v 5v 0ns 10us 10us 2ms 4ms  *input A
vb 4 0 pulse 0v 5v 0ns 10us 10us 4ms 8ms  *input B
*output at node 5
**********
mn1 5 3 0 0 nmod w=10u l=2u
mn2 5 4 0 0 nmod w=10u l=2u
mp1 2 3 1 1 pmod w=10u l=2u
mp2 5 4 2 1 pmod w=10u l=2u
**********
.model nmod nmos vto=1v kp=20u
.model pmod pmos vto=-1v kp=20u
.tran 0ns 8ms 10us 100us
.control
run
plot v(5) v(3) v(4)
.endc
.end
