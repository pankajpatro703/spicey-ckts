CMOS SR latch
*
*    Copyright (C) 2020, 2021 Pankajkumar Patro Licensed under the
*    Educational Community License, Version 2.0 (the "License"); you may
*    not use this file except in compliance with the License. You may
*    obtain a copy of the License at
*
*    http://www.osedu.org/licenses/ECL-2.0
*
*    Unless required by applicable law or agreed to in writing,
*    software distributed under the License is distributed on an "AS IS"
*    BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express
*    or implied. See the License for the specific language governing
*    permissions and limitations under the License.
*
***************************
* @Author: pankajpatro703 *
*  Released under ECL v2  *
***************************
vdd 1  0 dc    5v
*input S
vs  s  0 pulse 0v 5v 0ns 10us 10us 2ms 4ms
*input R
vr  r  0 pulse 0v 5v 0ns 10us 10us 1ms 2ms
*output at node Q, Q1
**********
* n-mos *
msn  q1  s   0   0  nmod w=10u l=2u
mrn  q   r   0   0  nmod w=10u l=2u
mqn  q1  q   0   0  nmod w=10u l=2u
mq1n q   q1  0   0  nmod w=10u l=2u
* p-mos *
msp  n1  s   1   1  pmod w=10u l=2u
mrp  n2  r   1   1  pmod w=10u l=2u
mqp  q1  q   n1  1  pmod w=10u l=2u
mq1p q   q1  n2  1  pmod w=10u l=2u
**********
.model nmod nmos vto=1v  kp=20u
.model pmod pmos vto=-1v kp=20u
.tran 1ns 4ms 10us 100us
.control
run
plot v(q) v(q1)
plot v(s) v(r)
.endc
.end
